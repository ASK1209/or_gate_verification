// Code your design here
module or_gate (
    input logic a,
    input logic b,
    output logic y
);
    assign y = a | b;
endmodule